//////
//ROM
/////

module Microstore_ROM (output reg[54:0] out, input [5:0] index);

initial begin

	//index =  6'b000001;
	
end

always @(index)

begin

	case(index)
		6'b000000:  out = 32'b00000000111100010000000000000000;
		6'b000001:  out = 32'b00010100011100000000000100111101;
		6'b000010:  out = 32'b11000000111100001000000000000000;
		6'b000011:  out = 32'b00000010110000000000000000000000;
		6'b000100:  out = 32'b00000100011100000000000000111101;
		6'b000101:  out = 32'b00000000111101000011000010100010;
		6'b000110:  out = 32'b00000100011100000000000000111101;
		6'b000111:  out = 32'b00000000111101000011000010111000;
		6'b001000:  out = 32'b00000000111100000000000000000000;
		6'b001001:  out = 32'b00000100011100000000000000111101;
		6'b001010:  out = 32'b00000000111101000110000010110100;
		6'b001011:  out = 32'b00000100011100000000000000111101;
		6'b001100:  out = 32'b00000100111100000000001100110010;
		6'b001101:  out = 32'b00000100011100000000000000111101;
		6'b001110:  out = 32'b00000100111100000000001100110100;
		6'b001111:  out = 32'b00000100111100000000001100110010;
		6'b010000:  out = 32'b00000100011100000000000000111101;
		6'b010001:  out = 32'b00000100111100000000001100110100;
		6'b010010:  out = 32'b00000100111100000000001100110010;
		6'b010011:  out = 32'b00000100111100000000001100110100;
		6'b010100:  out = 32'b00000000011100000000000010110010;
		6'b010101:  out = 32'b00000000011100000000000010110100;
		6'b010110:  out = 32'b00000100011100000000000000111101;
		6'b010111:  out = 32'b00000000111101000011000010110000;
		6'b011000:  out = 32'b00000100011100000000000000111101;
		6'b011001:  out = 32'b00000000111101000011000010110100;
		6'b011010:  out = 32'b00000000111101000011000010110010;
		6'b011011:  out = 32'b00000100011100000000000000111101;
		6'b011100:  out = 32'b00000000111101000011000010110100;
		6'b011101:  out = 32'b00000100011100000000000000111101;
		6'b011110:  out = 32'b00000000111100000000000000000000;
		6'b011111:  out = 32'b00000100111100000000001100110010;
		6'b100000:  out = 32'b00000100011100000000000000110101;
		6'b100001:  out = 32'b00000100111100000000001100110010;
		6'b100010:  out = 32'b00000100011100000000000000111101;
		6'b100011:  out = 32'b00000100111100000000001100110100;
		6'b100100:  out = 32'b00000100111100000000001100100010;
		6'b100101:  out = 32'b00000100111100000000001100110100;
		6'b100110:  out = 32'b00000000011100000000000010110010;
		6'b100111:  out = 32'b00000000011100000000000010110100;
		6'b101000:  out = 32'b00000100111100000010000100111101;
		6'b101001:  out = 32'b00000000111100000001010000100100;
		6'b101010:  out = 32'b00000000111100000001010000100100;
		6'b101011:  out = 32'b00100001111110000000000000110000;
		6'b101100:  out = 32'b00101100111110000000001100110000;

		6'
		
		
	endcase
end

endmodule
