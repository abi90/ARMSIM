module test_encoder;
wire [6:0] encOut;
reg [31:0]I;
encoder ec(encOut, I);
initial 
begin
#10 I <= 32'bxxxx01000x00xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0000100&&encOut), I, 7'b0000100,encOut);
#10 I <= 32'bxxxx01001x00xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0000110&&encOut), I, 7'b0000110,encOut);
#10 I <= 32'bxxxx01010x10xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0001000&&encOut), I, 7'b0001000,encOut);
#10 I <= 32'bxxxx01011x10xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0001010&&encOut), I, 7'b0001010,encOut);
#10 I <= 32'bxxxx01100x00xxxxxxxx00000000xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0001011&&encOut), I, 7'b0001011,encOut);
#10 I <= 32'bxxxx01101x00xxxxxxxx00000000xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0001101&&encOut), I, 7'b0001101,encOut);
#10 I <= 32'bxxxx01110x10xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0001111&&encOut), I, 7'b0001111,encOut);
#10 I <= 32'bxxxx01111x10xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0010001&&encOut), I, 7'b0010001,encOut);
#10 I <= 32'bxxxx01110x00xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0010010&&encOut), I, 7'b0010010,encOut);
#10 I <= 32'bxxxx01111x00xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0010011&&encOut), I, 7'b0010011,encOut);
#10 I <= 32'bxxxx01010x00xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0010100&&encOut), I, 7'b0010100,encOut);
#10 I <= 32'bxxxx01011x00xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0010101&&encOut), I, 7'b0010101,encOut);
#10 I <= 32'bxxxx01000x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0010110&&encOut), I, 7'b0010110,encOut);
#10 I <= 32'bxxxx01001x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0011000&&encOut), I, 7'b0011000,encOut);
#10 I <= 32'bxxxx01010x11xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0011010&&encOut), I, 7'b0011010,encOut);
#10 I <= 32'bxxxx01011x11xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0011100&&encOut), I, 7'b0011100,encOut);
#10 I <= 32'bxxxx01100x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0011101&&encOut), I, 7'b0011101,encOut);
#10 I <= 32'bxxxx01101x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0011111&&encOut), I, 7'b0011111,encOut);
#10 I <= 32'bxxxx01110x11xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0100001&&encOut), I, 7'b0100001,encOut);
#10 I <= 32'bxxxx01111x11xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0100011&&encOut), I, 7'b0100011,encOut);
#10 I <= 32'bxxxx01110x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0100100&&encOut), I, 7'b0100100,encOut);
#10 I <= 32'bxxxx01111x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0100101&&encOut), I, 7'b0100101,encOut);
#10 I <= 32'bxxxx01010x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0100110&&encOut), I, 7'b0100110,encOut);
#10 I <= 32'bxxxx01011x01xxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0100111&&encOut), I, 7'b0100111,encOut);
#10 I <= 32'bxxxx1011xxxxxxxx111xxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0101000&&encOut), I, 7'b0101000,encOut);
#10 I <= 32'bxxxx1010xxxxxxxx111xxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0101010&&encOut), I, 7'b0101010,encOut);
#10 I <= 32'bxxxx001xxxxxxxxxxxxxxxxxxxxxxxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0101011&&encOut), I, 7'b0101011,encOut);
#10 I <= 32'bxxxx000xxxxxxxxxxxxxxxxxxxx0xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0101100&&encOut), I, 7'b0101100,encOut);
#10 I <= 32'bxxxx00000100xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0101101&&encOut), I, 7'b0101101,encOut);
#10 I <= 32'bxxxx00001100xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0101111&&encOut), I, 7'b0101111,encOut);
#10 I <= 32'bxxxx00010110xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0110001&&encOut), I, 7'b0110001,encOut);
#10 I <= 32'bxxxx00011110xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0110011&&encOut), I, 7'b0110011,encOut);
#10 I <= 32'bxxxx00000000xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0110100&&encOut), I, 7'b0110100,encOut);
#10 I <= 32'bxxxx00001000xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0110110&&encOut), I, 7'b0110110,encOut);
#10 I <= 32'bxxxx00010010xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0111000&&encOut), I, 7'b0111000,encOut);
#10 I <= 32'bxxxx00011010xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0111010&&encOut), I, 7'b0111010,encOut);
#10 I <= 32'bxxxx00010000xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0111011&&encOut), I, 7'b0111011,encOut);
#10 I <= 32'bxxxx00011000xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0111100&&encOut), I, 7'b0111100,encOut);
#10 I <= 32'bxxxx00010100xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0111101&&encOut), I, 7'b0111101,encOut);
#10 I <= 32'bxxxx00011100xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0111110&&encOut), I, 7'b0111110,encOut);
#10 I <= 32'bxxxx00000101xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (0111111&&encOut), I, 7'b0111111,encOut);
#10 I <= 32'bxxxx00001101xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1000001&&encOut), I, 7'b1000001,encOut);
#10 I <= 32'bxxxx00010111xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1000011&&encOut), I, 7'b1000011,encOut);
#10 I <= 32'bxxxx00011111xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1000101&&encOut), I, 7'b1000101,encOut);
#10 I <= 32'bxxxx00000001xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1000110&&encOut), I, 7'b1000110,encOut);
#10 I <= 32'bxxxx00001001xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1001000&&encOut), I, 7'b1001000,encOut);
#10 I <= 32'bxxxx00010011xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1001010&&encOut), I, 7'b1001010,encOut);
#10 I <= 32'bxxxx00011011xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1001100&&encOut), I, 7'b1001100,encOut);
#10 I <= 32'bxxxx00010001xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1001101&&encOut), I, 7'b1001101,encOut);
#10 I <= 32'bxxxx00011001xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1001110&&encOut), I, 7'b1001110,encOut);
#10 I <= 32'bxxxx00010101xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1001111&&encOut), I, 7'b1001111,encOut);
#10 I <= 32'bxxxx00011101xxxxxxxxxxxx1xx1xxxx;
#10 $display("Test Result=%b I=%b Expected=%b Result=%b", (1010000&&encOut), I, 7'b1010000,encOut);
end																	
endmodule